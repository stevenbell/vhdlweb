module add1 (input logic[7:0] operand,
             output logic[7:0] result);

    assign result = operand + 1;

endmodule


